package processor_test_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"

  import processor_agent_pkg::*;
  import processor_env_pkg::*;

  `include "processor_sequence.sv"
  `include "processor_test.sv"
endpackage