package processor_env_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"

  import processor_agent_pkg::*;

  `include "processor_scoreboard.sv"
  `include "processor_subscriber.sv"
  `include "processor_env.sv"
endpackage