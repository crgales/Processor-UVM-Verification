package processor_agent_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"
  
  `include "processor_transaction.sv"
  `include "processor_driver.sv"
  `include "processor_monitor.sv"
  `include "processor_agent.sv"
endpackage
  
